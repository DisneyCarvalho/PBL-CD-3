module pulse(Clock, Level, Pulse);
	input Clock, Level;
	output Pulse;
	
	reg [1:0] state, nextstate;
	
	parameter S0 =2'b00;
	parameter S1 =2'b01;
	parameter S2 =2'b10;
	

	
	// state register
	always @ ( posedge Clock)	
		state <= nextstate ;
		
	// next state logic
	always @ (*)
		case ( state )
			S0 : if ( Level ) nextstate <= S1 ;
			else nextstate <= S0 ;
			S1 : if ( Level ) nextstate <= S2 ;
			else nextstate <= S0 ;
			S2 : if ( Level ) nextstate <= S2 ;
			else nextstate <= S0 ;
			default : nextstate <= S0 ;
			
		endcase
		
	// output logic
	assign Pulse = ( state == S1 ) ;
	endmodule